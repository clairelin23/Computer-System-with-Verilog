`timescale 1ns/1ps

module mux_1b_tb;

/*
//output list
wire Y;
//input list
reg I0, I1, S;

MUX1_2x1 inst1(Y,I0, I1, S);

initial
begin
I0=0; I1=1; S =0;
#5 I0=0; I1=1; S =1;
#5 I0=1; I1=0; S =0;
#5 I0=1; I1=0; S =1;
end
endmodule

wire [31:0] Y;
//input list
reg [31:0] I0, I1;
reg  S;

MUX32_2x1 inst1(Y, I0, I1, S);

initial
begin
I0=0; I1=10; S =0;
#5 I0=5; I1=100; S =1;
#5 I0=5; I1=100; S =0;
#5 I0=15; I1=8; S =1;
end
endmodule


//input list
reg [31:0] I0, I1, I2, I3;
reg [1:0] S;
wire [31:0] Y;

MUX32_4x1 inst1 (Y, I0, I1, I2, I3, S);


initial
begin
I0=0; I1=0; I2 = 0; I3 = 0; S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; S =1;
#5 I0=5; I1=100; I2 = 30; I3 = 40; S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; S =2;
#5 I0=5; I1=100; I2 = 30; I3 = 40; S =3;
#5;
end
endmodule


//input list
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7;
reg [2:0] S;
wire [31:0] Y;

// 32-bit 8x1 mux
MUX32_8x1 inst1(Y, I0, I1, I2, I3, I4, I5, I6, I7, S);


initial
begin
I0=0; I1=0; I2 = 0; I3 = 0; I4 =0; I5 = 9; I6= 8; I7=1; S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; S =1;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1;S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1;S =2;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; S =3;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; S =4;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; S =5;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; S =6;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; S =7;
#5;
end
endmodule


// 32-bit 16x1 mux
//input list
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7,I8, I9, I10, I11, I12, I13, I14, I15;
reg [3:0] S;
wire [31:0] Y;

MUX32_16x1 inst1 (Y, I0, I1, I2, I3, I4, I5, I6, I7,
                     I8, I9, I10, I11, I12, I13, I14, I15, S);


initial
begin
I0=0; I1=0; I2 = 0; I3 = 0; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 0; I9=0; I10=0; I11=0; I12=0; I13=0; I14=3; I15=3; S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; S =1;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =2;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =3;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =4;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =5;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =6;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =7;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =8;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =9;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =10;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =11;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =12;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =13;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =14;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;S =15;
#5;
end
*/

// output list
wire [31:0] Y;
//input list
reg [31:0] I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15;
reg [31:0] I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31;
reg [4:0] S;
 MUX32_32x1 inst11(Y, I0, I1, I2, I3, I4, I5, I6, I7,
                     I8, I9, I10, I11, I12, I13, I14, I15,
                     I16, I17, I18, I19, I20, I21, I22, I23,
                     I24, I25, I26, I27, I28, I29, I30, I31, S);


initial
begin
I0=0; I1=0; I2 = 0; I3 = 0; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 0; I9=0; I10=0; I11=0; I12=0; I13=0; I14=3; I15=3; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44; S = 0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44; S =1;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =0;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =2;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =3;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =4;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;  I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =5;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =6;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;  I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =7;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;  I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =8;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;  I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =9;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;  I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =10;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =11;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =12;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28;  I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =13;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =14;
#5 I0=5; I1=100; I2 = 30; I3 = 40; I4 =0; I5 = 9; I6= 8; I7=1; I8 = 21; I9=22; I10=23; I11=24; I12=25; I13=26; I14=27; I15=28; I16 = 29; I17 =30; I18 = 31; I19= 32; I20=33; I21 = 34; I22=35; I23=36; I24=37; I25=38; I26=39; I27=40; I28=41 ;I29 =42; I30 = 43; I31 = 44;S =31;
#5;
end
endmodule


